package ALU_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"

    `include "ALU_Sequence_Item.sv"
    `include "ALU_Sequence.sv"
    `include "ALU_Sequencer.sv"
    `include "ALU_Driver.sv"
    `include "ALU_monitor.sv"
    `include "ALU_Coverage_Collector.sv"
    `include "ALU_Scoreboard.sv"
    `include "ALU_Agent.sv"
    `include "ALU_Env.sv"
    `include "Test.sv"
endpackage: ALU_pkg
